`include "test_ldi.vh"
`include "test_in.vh"
`include "test_out.vh"
